`timescale 1ns/100ps

`include "define_drive_circuit_inst_decoder.v"

module drive_circuit_inst_decoder_tb();
// TODO
endmodule
